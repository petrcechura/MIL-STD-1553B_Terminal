library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

--Model is divided into two parts - Synchronize detector and Manchester decoder; first part is used for detection of synchronize waveform which stands
--for 3 bits. Detection is realized by state machine and timer; when a pos or neg input occurs, timer runs until 3/2 period (see Word Formats),
--then state is changed and opposite value is required. Whenever anything unexpected happens, state returns to default. Whenever a full synchronize waveform is detected, 
--data are sent to the second part, but only for 17 bit periods; after that time, state is returned to the default.
--Second part is free of any state machine and just gets log. value in every 3/4 period of data; output is then decoded signal.

--Sync type carries information how synchronization begins (data word begins with neg waveform, command with pos waveform)

entity ManchesterDecoder is
    -- for frequency 1 MHz
    port (
        clk   : in std_logic;
        reset : in std_logic;
        in_positive, in_negative : in std_logic;
        data_out : out std_logic;
        RX_done : out std_logic;
        state_out : out std_logic_vector(2 downto 0)
    );
end entity;



architecture rtl of ManchesterDecoder is
    -- SYNCHRONIZE DETECTOR --
    type t_state is (s_default, --default state, terminal is waiting for signal
                     s_logic_one1, --
                     s_logic_one2,
                     s_logic_one3, 
                     s_logic_two1, 
                     s_logic_two2,
                     s_logic_two3, 
                     s_synchronize); -- stands for 17 manchester bit periods (measured just by time and known frequency); then goes to default
    signal state_q, state_d : t_state;

    --timer for sync sample
    signal sync_timer_en : std_logic;
    signal sync_timer_d, sync_timer_q : unsigned(4 downto 0);
    signal sync_timer_max : std_logic;

    -- MANCHESTER DECODER --
    --timer for data sample
    signal manchester_timer_en : std_logic;
    signal manchester_timer_d, manchester_timer_q : unsigned(4 downto 0);
    signal manchester_timer_sample : std_logic;

    --counter for data count
    signal data_counter_en : std_logic;
    signal data_counter_d, data_counter_q : unsigned(3 downto 0); -- counts to 16 (16-bit word)
    signal data_counter_max : std_logic;
    --data register
    signal decoded_data : unsigned(3 downto 0);




    
begin

    --*** SYNCHRONIZE DETECTOR ***--

    -- MAIN STATE MACHINE
    --seq part
    process (clk)
    begin
        if reset='1' then
            state_q <= s_default;
        elsif rising_edge(clk) then
            state_q <= state_d;
        end if;
    end process;

    --comb part
    process (state_q)
    begin
        case state_q is 
            when s_default =>
                sync_timer_en <= '0';
                manchester_timer_en <= '0';

                if in_positive= '1' and in_negative='0' then
                    state_d <= s_logic_one1;
                elsif in_negative = '1' and in_positive = '0' then
                    state_d <= s_logic_two1;
                else
                    state_d <= s_default;
                end if;
            when s_logic_one1 =>
                sync_timer_en <= '1';
                manchester_timer_en <= '0';

                if sync_timer_max='1' then
                    state_d <= s_logic_one2;
                elsif in_positive='1' and in_negative='0' then
                    state_d <= s_logic_one1;
                else
                    state_d <= s_default;
                end if;

            when s_logic_one2 =>
                sync_timer_en <= '1';
                manchester_timer_en <= '0';

                if sync_timer_max='1' then
                    state_d <= s_logic_one3;
                else
                    state_d <= s_logic_one2;
                end if;

            when s_logic_one3 =>
                sync_timer_en <= '1';
                manchester_timer_en <= '0';

                if sync_timer_max='1' then
                    state_d <= s_synchronize;
                elsif in_positive='0' and in_negative='1' then
                    state_d <= s_logic_one3;
                else
                    state_d <= s_default;
                end if;

            when s_logic_two1 =>
                sync_timer_en <= '1';
                manchester_timer_en <= '0';

                if sync_timer_max='1' then
                    state_d <= s_logic_two2;
                elsif in_positive='0' and in_negative='1' then
                    state_d <= s_logic_two1;
                else
                    state_d <= s_default;
                end if;
            when s_logic_two2 =>
                sync_timer_en <= '1';
                manchester_timer_en <= '0';

                if sync_timer_max='1' then
                    state_d <= s_logic_two3;
                else
                    state_d <= s_logic_two2;
                end if;
            when s_logic_two3 =>
                sync_timer_en <= '1';
                manchester_timer_en <= '0';

                if sync_timer_max='1' then
                    state_d <= s_synchronize;
                elsif in_positive='1' and in_negative='0' then
                    state_d <= s_logic_two3;
                else
                    state_d <= s_default;
                end if;

            when s_synchronize =>
                sync_timer_en <= '0';
                manchester_timer_en <= '1';


        end case;
    end process;

    -- SYNC TIMER SAMPLE
    --seq part
    process (clk)
    begin
        if reset='1' then
            sync_timer_q <= (others => '0'); 
        elsif rising_edge(clk) then
            sync_timer_q <= sync_timer_d;
        end if;
    end process;

    -- comb part
    process (sync_timer_q)
    begin
        if sync_timer_en='1' then
            sync_timer_d <= sync_timer_q+1;
        else
            sync_timer_d <= (others => '0');
        end if; 

        if sync_timer_q = (others => '1') then
            sync_timer_max <= '1';
        end if;

    end process;

    --- *** MANCHESTER SAMPLE *** ---

    -- MANCHESTER TIMER SAMPLE
    --seq part
    process (clk)
    begin
        if reset='1' then
            manchester_timer_q <= (others => '0'); 
        elsif rising_edge(clk) then
            manchester_timer_q <= manchester_timer_d;
        end if;
    end process;

    --comb part
    process (manchester_timer_q)
    begin
        if manchester_timer_en='1' then
            manchester_timer_d <= manchester_timer_q + 1;
        else
            manchester_timer_d <= (others => '0'); 
        end if;

        if manchester_timer_q=24 then
            manchester_timer_sample <= '1';
        else
            manchester_timer_sample <= '0';
        end if;

    end process;

    -- DATA REGISTER
    process (clk)
    begin
        if rising_edge(clk) then
            
        end if;
    end process;





end architecture;
